/*
 * Copyright 2017 IBM Corporation
 * Licensed to the Apache Software Foundation (ASF) under one
 * or more contributor license agreements.  See the NOTICE file
 * distributed with this work for additional information
 * regarding copyright ownership.  The ASF licenses this file
 * to you under the Apache License, Version 2.0 (the
 * "License"); you may not use this file except in compliance
 * with the License.  You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * Author: Andrew K Martin akmartin@us.ibm.com
 */
 
module base_vlat_rst #
  (   parameter width=1
   )
   (
    input 	       clk,
    input 	       reset,
    input [width-1:0]  din,
    input [width-1:0]  rstv,
    output [width-1:0] q
    );
   

   reg [width-1:0]    q_int;

   always@(posedge clk or posedge reset)
     if (reset) q_int <= rstv;
     else q_int <= din;
   assign q = q_int;
   
endmodule // base_vlat


   
  

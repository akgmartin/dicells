/*
 * Copyright 2017 IBM Corporation
 * Licensed to the Apache Software Foundation (ASF) under one
 * or more contributor license agreements.  See the NOTICE file
 * distributed with this work for additional information
 * regarding copyright ownership.  The ASF licenses this file
 * to you under the Apache License, Version 2.0 (the
 * "License"); you may not use this file except in compliance
 * with the License.  You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * Author: Andrew K Martin akmartin@us.ibm.com
 */
 
module base_pridemux#
  (   
      parameter ways = 2,
      parameter width = 1
      )
   (
    input 	       i_v,
    output 	       i_r,
    output [0:ways-1]  o_v,
    input [0:ways-1]   o_r
   );

   wire [0:ways-1]     s1_r;
   
   base_priarb#(.ways(ways)) iarb
     (.i_v(o_r), .i_r(o_v),
      .o_v(s1_r), .o_r(i_v)
      );
   assign i_r = | s1_r;
   
endmodule // base_pri_arb

		     
